module main();


endmodule